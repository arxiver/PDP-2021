library ieee;
use ieee.std_logic_1164.ALL;
use ieee.numeric_std.all;

entity RomEnt is
    port(
            Clk : in std_logic;
            Address : in std_logic_vector(7 downto 0);
            Output : out std_logic_vector(24 downto 0)
        );
end entity;

architecture RomArc of RomEnt is

type RomType is array(0 to 256) of std_logic_vector(24 downto 0);   -- 40
signal Rom : RomType:=
(
    --              F8           F1      F2      F3      F4      F5      F6      F7
    0   =>	"00000001" &	"001" &	"011" &	"01" &	"00" &	"01" &	"01" &	"000",
    1   =>	"00000010" &	"011" &	"001" &	"00" &	"01" &	"00" &	"00" &	"000",
    2   =>	"00000011" &	"010" &	"010" &	"00" &	"00" &	"00" &	"00" &	"000",
    3   =>	"11111111" &    "000" &	"000" &	"00" &	"00" &	"00" &	"00" &	"101",
    40  =>      "00101001" &	"111" &	"011" &	"00" &	"00" &	"11" &	"00" &	"000",
    41  =>	"00000000" &	"011" &	"001" &	"00" &	"00" &	"00" &	"00" &	"000",
    48  =>      "00000000" &    "000" &"000" &	"00" &	"00" &	"00" &	"00" &	"000",
    65  =>	"01111000" &	"100" &	"000" &	"00" &	"10" &	"00" &	"00" &	"001",
    73  =>	"01110110" &    "100" &	"000" &	"01" &	"00" &	"00" &	"01" &	"010", -- base address 166
    81 =>	"01010010" &    "100" &	"011" &	"01" &	"01" &	"01" &	"01" &	"000",
    82  =>	"01110110" &    "011" &	"100" &	"00" &	"00" &	"00" &	"00" &	"010", -- base address 166
    97  =>	"01100010" &	"100" &	"011" &	"00" &	"01" &	"10" &	"00" &	"000",
    98  =>	"01110110" &    "011" &	"100" &	"01" &	"00" &	"00" &	"01" &	"010", -- base address 166
    113 =>	"01110010" &	"001" &	"011" &	"01" &	"01" &	"01" &	"01" &	"000",
    114 =>	"01110011" &	"011" &	"001" &	"00" &	"00" &	"00" &	"00" &	"000",
    115 =>	"01110100" &	"010" &	"000" &	"00" &	"01" &	"00" &	"00" &	"000",
    116 =>	"01110101" &	"100" &	"011" &	"00" &	"00" &	"00" &	"00" &	"000",
    117 =>	"01110110" &    "011" &	"000" &	"01" &	"00" &	"00" &	"01" &	"010", -- base address 166
    118 =>	"01110111" &	"010" &	"000" &	"01" &	"00" &	"00" &	"01" &	"000",
    119 =>	"01111000" &	"010" &	"000" &	"00" &	"10" &	"00" &	"00" &	"001",
    -- 170 =>	"GO TO BETA" &							-	,
    129 =>	"10111000" &	"101" &	"000" &	"00" &	"01" &	"00" &	"00" &	"000",
    137 =>	"10110111" &    "101" &	"000" &	"01" &	"00" &	"00" &	"01" &	"000", -- base address 266
    145 =>	"10010010" &	"101" &	"011" &	"01" &	"01" &	"01" &	"01" &	"000",
    146 =>	"10110110" &    "011" &	"101" &	"00" &	"00" &	"00" &	"00" &	"011", -- base address 266
    161 =>	"10100010" &	"101" &	"011" &	"00" &	"01" &	"10" &	"00" &	"000",
    162 =>	"10110110" &    "011" &	"101" &	"01" &	"00" &	"00" &	"01" &	"011", -- base address 266
    177 =>	"10110010" &	"001" &	"011" &	"01" &	"01" &	"01" &	"01" &	"000",
    178 =>	"10110011" &	"011" &	"001" &	"00" &	"00" &	"00" &	"00" &	"000",
    179 =>	"10110100" &	"010" &	"000" &	"00" &	"01" &	"00" &	"00" &	"000",
    180 =>	"10110101" &	"101" &	"011" &	"00" &	"00" &	"00" &	"00" &	"000",
    181 =>	"10110110" &    "011" &	"000" &	"01" &	"00" &	"00" &	"01" &	"011", -- base address 266
    182 =>	"10110111" &	"010" &	"000" &	"01" &	"00" &	"00" &	"01" &	"000",
    183 =>	"10111000" &	"010" &	"000" &	"00" &	"01" &	"00" &	"00" &	"000",
    184 =>	"10111010" &    "110" &	"011" &	"00" &	"00" &	"11" &	"00" &	"100", -- base address 271
    186 =>	"00000000" &	"011" &	"000" &	"10" &	"00" &	"00" &	"10" &	"000",
    187 =>	"00000000" &	"011" &	"101" &	"00" &	"00" &	"00" &	"00" &	"000",
    188 =>	"00000000" &	"000" &	"000" &	"00" &	"00" &	"00" &	"00" &	"000",
    others => "0000000000000000000000000"
);


begin
    process(Clk) is
    begin
        if rising_edge(Clk) then
            Output <= Rom(to_integer(unsigned((Address))));
        end if;
    end process;
end RomArc;